`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:05:02 10/31/2020 
// Design Name: 
// Module Name:    Procesador 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Procesador(
    input [31:0] Data_in,
    input Clk,
    input Reset,
    output [5:0] Address,
    output [31:0] Data_out,
    output We
    );


endmodule
